//a Note: created by CDL 1.4 - do not hand edit without recognizing it will be out of sync with the source
// Output mode 0 (VMOD=1, standard verilog=0)
// Verilog option comb reg suffix '__var'
// Verilog option include_displays 0
// Verilog option include_assertions 1
// Verilog option sv_assertions 0
// Verilog option assert delay string '<NULL>'
// Verilog option include_coverage 0
// Verilog option clock_gate_module_instance_type 'banana'
// Verilog option clock_gate_module_instance_extra_ports ''
// Verilog option use_always_at_star 1
// Verilog option clocks_must_have_enables 1

//a Module led_ws2812_chain
    //   
    //   A chain of any length of Neopixel LEDs can be driven by this module
    //   
    //   The interface is a request/data interface; this module presents a
    //   @a ready request to the client, which then presents a valid 24-bit
    //   RGB data value. When the module takes the data it removes its
    //   @a ready request. The client keeps supplying data in response to the
    //   @a ready requests.
    //    
    //   To terminate the chain the client supplies data with a @a last
    //   indication asserted.
    //   
    //   To ease implementation of the client, the request includes a
    //   @a first indicator and an @a led_number indicator - effectively a
    //   client can read a register file based on @a led_number and drive
    //   @a valid when the data is valid, and @a last if led_number matches
    //   the end of the register file.
    //   
    //   This module copes with all of the requirements of the Neopixel
    //   chain, and it takes a constant clock input. To provide the correct
    //   frequency of data pin toggling to the Neopixels a clock divider
    //   value must be supplied, with the approximate number of clock ticks
    //   that make up 400ns (ideally 408ns).
    //   
    //   The Neopixel WS2812 LED chains use a serial data stream with encoded
    //   clock to provide data to the LEDs.
    //   
    //   If the LED chain data is held low for >50us then the stream performs a
    //   'load to LEDs' - this transfers the serial data already loaded in to
    //   the LEDs to the actual LED drivers themselves.
    //   
    //   Before loading the LEDs the chain should be fed data.  The data is fed
    //   using a high/low data pulse per bit. The ratio high/low provides the
    //   data bit value.
    //   
    //   A high/low of 1:2 provids a zero bit; a high/low of 1:2 provides a one
    //   bit. The total bit time should be 1.25us.  Hence this logic requires a
    //   1.25/3us, or roughly 400ns clock generator. This is performed using a
    //   clock divider and a user-supplied divide value, which will depend on
    //   the input clock frequency. For example, if the input clock frequency
    //   is 50MHz, which is a period of 20ns, then the divider should be set to
    //   20.
    //   
    //   The data is provided to the LEDs green, red then blue, most
    //   significant bit first, with 8 bits for each component.
    //   
    //   The logic uses a simple state machine; when it is idle it will have no
    //   data in hand, and need data to feed in to the LED stream. At this
    //   point it requests a valid first LED data. When valid data is received
    //   into a buffer the state machine transitions to the data-in-hand state;
    //   it remains there until the data transmitter takes the data, when it
    //   either requests more data (as per idle), or if the last LED data was
    //   provided by the client, it moves to requests an LED load, and it waits
    //   in loading state until that completes. At this point it transitions
    //   back to idle, and the process restarts.
    //   
    //   When there is valid LED data in the internal buffer the data
    //   transmitter can start; the data is transferred to the shift register,
    //   and it is driven out by the data transmitter to the LED chain one bit
    //   at a time.
    //   
    //   
module led_ws2812_chain
(
    clk,
    clk__enable,

    led_data__valid,
    led_data__last,
    led_data__red,
    led_data__green,
    led_data__blue,
    divider_400ns,
    reset_n,

    led_chain,
    led_request__ready,
    led_request__first,
    led_request__led_number
);

    //b Clocks
        //   System clock - not the pin clock, which is derived from this
    input clk;
    input clk__enable;

    //b Inputs
        //   LED data, for the requested led
    input led_data__valid;
    input led_data__last;
    input [7:0]led_data__red;
    input [7:0]led_data__green;
    input [7:0]led_data__blue;
        //   clock divider value to provide for generating a pulse every 400ns based on clk
    input [7:0]divider_400ns;
        //   Active low reset
    input reset_n;

    //b Outputs
        //   Data pin for LED chain, modulated by this module to drive LED settings
    output led_chain;
        //   LED data request, to get data from the next LED to light
    output led_request__ready;
    output led_request__first;
    output [7:0]led_request__led_number;

// output components here

    //b Output combinatorials
        //   Data pin for LED chain, modulated by this module to drive LED settings
    reg led_chain;
        //   LED data request, to get data from the next LED to light
    reg led_request__ready;
    reg led_request__first;
    reg [7:0]led_request__led_number;

    //b Output nets

    //b Internal and output registers
        //   Modulator (data_chain) state
    reg [7:0]data_chain_state__divider;
    reg data_chain_state__active;
    reg data_chain_state__sr__valid;
    reg [2:0]data_chain_state__sr__value;
    reg [1:0]data_chain_state__value_number;
    reg data_chain_state__output_data;
        //   Transmitter state, the state of the internal transmit state machine
    reg [2:0]data_transmitter_state__fsm_state;
    reg data_transmitter_state__shift_register__valid;
    reg data_transmitter_state__shift_register__last;
    reg [7:0]data_transmitter_state__shift_register__red;
    reg [7:0]data_transmitter_state__shift_register__green;
    reg [7:0]data_transmitter_state__shift_register__blue;
    reg [5:0]data_transmitter_state__counter;
        //   Data state, the state of the interface to the client
    reg [1:0]data_state__fsm_state;
    reg [7:0]data_state__led_number;
    reg data_state__buffer__valid;
    reg data_state__buffer__last;
    reg [7:0]data_state__buffer__red;
    reg [7:0]data_state__buffer__green;
    reg [7:0]data_state__buffer__blue;
    reg data_state__load_leds;

    //b Internal combinatorials
        //   Combinatorial decode of modulator state
    reg data_chain_combs__clk_enable;
    reg data_chain_combs__taking_transmitter_data;
        //   Combinatorial decode of the transmitter state
    reg data_transmitter_combs__loading_leds;
    reg data_transmitter_combs__taking_data;
    reg data_transmitter_combs__needs_data;
    reg data_transmitter_combs__idle_transmitter;
    reg data_transmitter_combs__selected_data;
    reg data_transmitter_combs__load_leds;
    reg data_transmitter_combs__drive_bits__valid;
    reg [2:0]data_transmitter_combs__drive_bits__value;
    reg data_transmitter_combs__counter_expired;

    //b Internal nets

    //b Clock gating module instances
    //b Module instances
    //b data_state_machine_logic__comb combinatorial process
        //   
        //       The data state machine is a simple interface to the led request
        //       and led_data, feeding the data transmitter shift register when it
        //       can.
        //   
        //       It has a data_buffer that it stores incoming led data in, and it
        //       feeds this to the data transmitter shift register when permitted,
        //       invalidating the data buffer.
        //   
        //       If the transmitter takes a @a last data then the state machine will
        //       then request that the transmitter 'load the leds'; this request
        //       will, of course, have to wait for the completion of the current
        //       shift register contents (the last LED), and then the correct 50us
        //       of data will presumably be transmitted. During this time the data
        //       state machine can be requesting the next set of data to transmit.
        //       So that the next LED data does not get too stale, the request
        //       should occur towards the end of the 50us of 'load led' - which it
        //       will do, as the transmitter state machine indicates that the LEDS
        //       are being loaded in the last microsecond of so of the 50us of
        //       'load led' time.
        //       
    always @ ( * )//data_state_machine_logic__comb
    begin: data_state_machine_logic__comb_code
    reg led_request__ready__var;
    reg led_request__first__var;
        led_request__ready__var = 1'h0;
        led_request__first__var = 1'h0;
        led_request__led_number = data_state__led_number;
        case (data_state__fsm_state) //synopsys parallel_case
        2'h0: // req 1
            begin
            led_request__ready__var = 1'h1;
            led_request__first__var = 1'h1;
            end
        2'h1: // req 1
            begin
            led_request__ready__var = 1'h1;
            led_request__first__var = 1'h0;
            end
        2'h2: // req 1
            begin
            end
        2'h3: // req 1
            begin
            end
    //synopsys  translate_off
    //pragma coverage off
        default:
            begin
                if (1)
                begin
                    $display("%t *********CDL ASSERTION FAILURE:led_ws2812_chain:data_state_machine_logic: Full switch statement did not cover all values", $time);
                end
            end
    //pragma coverage on
    //synopsys  translate_on
        endcase
        led_request__ready = led_request__ready__var;
        led_request__first = led_request__first__var;
    end //always

    //b data_state_machine_logic__posedge_clk_active_low_reset_n clock process
        //   
        //       The data state machine is a simple interface to the led request
        //       and led_data, feeding the data transmitter shift register when it
        //       can.
        //   
        //       It has a data_buffer that it stores incoming led data in, and it
        //       feeds this to the data transmitter shift register when permitted,
        //       invalidating the data buffer.
        //   
        //       If the transmitter takes a @a last data then the state machine will
        //       then request that the transmitter 'load the leds'; this request
        //       will, of course, have to wait for the completion of the current
        //       shift register contents (the last LED), and then the correct 50us
        //       of data will presumably be transmitted. During this time the data
        //       state machine can be requesting the next set of data to transmit.
        //       So that the next LED data does not get too stale, the request
        //       should occur towards the end of the 50us of 'load led' - which it
        //       will do, as the transmitter state machine indicates that the LEDS
        //       are being loaded in the last microsecond of so of the 50us of
        //       'load led' time.
        //       
    always @( posedge clk or negedge reset_n)
    begin : data_state_machine_logic__posedge_clk_active_low_reset_n__code
        if (reset_n==1'b0)
        begin
            data_state__fsm_state <= 2'h0;
            data_state__fsm_state <= 2'h0;
            data_state__led_number <= 8'h0;
            data_state__load_leds <= 1'h0;
            data_state__buffer__valid <= 1'h0;
            data_state__buffer__last <= 1'h0;
            data_state__buffer__red <= 8'h0;
            data_state__buffer__green <= 8'h0;
            data_state__buffer__blue <= 8'h0;
        end
        else if (clk__enable)
        begin
            case (data_state__fsm_state) //synopsys parallel_case
            2'h0: // req 1
                begin
                if ((led_data__valid!=1'h0))
                begin
                    data_state__fsm_state <= 2'h2;
                end //if
                end
            2'h1: // req 1
                begin
                if ((led_data__valid!=1'h0))
                begin
                    data_state__fsm_state <= 2'h2;
                end //if
                end
            2'h2: // req 1
                begin
                if (!(data_state__buffer__valid!=1'h0))
                begin
                    data_state__led_number <= (data_state__led_number+8'h1);
                    data_state__fsm_state <= 2'h1;
                    if ((data_state__buffer__last!=1'h0))
                    begin
                        data_state__fsm_state <= 2'h3;
                    end //if
                end //if
                end
            2'h3: // req 1
                begin
                data_state__load_leds <= 1'h1;
                if ((data_transmitter_combs__loading_leds!=1'h0))
                begin
                    data_state__load_leds <= 1'h0;
                    data_state__led_number <= 8'h0;
                    data_state__fsm_state <= 2'h0;
                end //if
                end
    //synopsys  translate_off
    //pragma coverage off
            default:
                begin
                    if (1)
                    begin
                        $display("%t *********CDL ASSERTION FAILURE:led_ws2812_chain:data_state_machine_logic: Full switch statement did not cover all values", $time);
                    end
                end
    //pragma coverage on
    //synopsys  translate_on
            endcase
            if (((led_request__ready!=1'h0)&&(led_data__valid!=1'h0)))
            begin
                data_state__buffer__valid <= led_data__valid;
                data_state__buffer__last <= led_data__last;
                data_state__buffer__red <= led_data__red;
                data_state__buffer__green <= led_data__green;
                data_state__buffer__blue <= led_data__blue;
            end //if
            if ((data_transmitter_combs__taking_data!=1'h0))
            begin
                data_state__buffer__valid <= 1'h0;
            end //if
        end //if
    end //always

    //b data_transmitter_logic__comb combinatorial process
        //   
        //       The data transmitter is responsible for reading data bits to the
        //       Neopixel data chain driver (modulator).
        //   
        //       It maintains a shift register (with separate @a red, @a green and @a blue
        //       components), with a @a valid bit.
        //   
        //       Data is loaded into the shift register when it is not valid. The
        //       transmitter then shifts straight in to asking the drive chain to
        //       output @a green[7]. It shifts the @a green bits up every time the
        //       drive chain takes a bit, and after 8 bits it moves to the @a red,
        //       and then the @a blue. At the end of the @a blue it invalidates the
        //       shift register.
        //   
        //       The shift register should be filled quickly enough for the data
        //       chain to not miss a beat, if further LED data is to be driven.
        //   
        //       Instead of driving out a shift register the state machine may be
        //       requested to drive out a 'load leds' value. This is 50us of 'low'
        //       on the output, which is achieved here by roughly 40 sets of drives
        //       of '0' for 1.25us each.
        //       
    always @ ( * )//data_transmitter_logic__comb
    begin: data_transmitter_logic__comb_code
    reg data_transmitter_combs__idle_transmitter__var;
    reg data_transmitter_combs__selected_data__var;
    reg data_transmitter_combs__load_leds__var;
    reg data_transmitter_combs__drive_bits__valid__var;
    reg [2:0]data_transmitter_combs__drive_bits__value__var;
    reg data_transmitter_combs__loading_leds__var;
        data_transmitter_combs__needs_data = !(data_transmitter_state__shift_register__valid!=1'h0);
        data_transmitter_combs__taking_data = ((data_state__buffer__valid!=1'h0)&&(data_transmitter_combs__needs_data!=1'h0));
        data_transmitter_combs__counter_expired = (data_transmitter_state__counter==6'h0);
        data_transmitter_combs__idle_transmitter__var = 1'h0;
        data_transmitter_combs__selected_data__var = 1'h0;
        data_transmitter_combs__load_leds__var = 1'h0;
        case (data_transmitter_state__fsm_state) //synopsys parallel_case
        3'h0: // req 1
            begin
            data_transmitter_combs__idle_transmitter__var = 1'h1;
            end
        3'h1: // req 1
            begin
            data_transmitter_combs__idle_transmitter__var = 1'h0;
            data_transmitter_combs__selected_data__var = data_transmitter_state__shift_register__green[7];
            end
        3'h2: // req 1
            begin
            data_transmitter_combs__idle_transmitter__var = 1'h0;
            data_transmitter_combs__selected_data__var = data_transmitter_state__shift_register__red[7];
            end
        3'h3: // req 1
            begin
            data_transmitter_combs__idle_transmitter__var = 1'h0;
            data_transmitter_combs__selected_data__var = data_transmitter_state__shift_register__blue[7];
            end
        3'h4: // req 1
            begin
            data_transmitter_combs__load_leds__var = 1'h1;
            end
    //synopsys  translate_off
    //pragma coverage off
        default:
            begin
                if (1)
                begin
                    $display("%t *********CDL ASSERTION FAILURE:led_ws2812_chain:data_transmitter_logic: Full switch statement did not cover all values", $time);
                end
            end
    //pragma coverage on
    //synopsys  translate_on
        endcase
        data_transmitter_combs__drive_bits__valid__var = 1'h0;
        data_transmitter_combs__drive_bits__value__var = 3'h0;
        if ((data_transmitter_combs__load_leds__var!=1'h0))
        begin
            data_transmitter_combs__drive_bits__valid__var = 1'h1;
            data_transmitter_combs__drive_bits__value__var = 3'h0;
        end //if
        else
        
        begin
            if (!(data_transmitter_combs__idle_transmitter__var!=1'h0))
            begin
                data_transmitter_combs__drive_bits__valid__var = 1'h1;
                data_transmitter_combs__drive_bits__value__var = {{1'h0,data_transmitter_combs__selected_data__var},1'h1};
            end //if
        end //else
        data_transmitter_combs__loading_leds__var = 1'h0;
        case (data_transmitter_state__fsm_state) //synopsys parallel_case
        3'h0: // req 1
            begin
            end
        3'h1: // req 1
            begin
            end
        3'h2: // req 1
            begin
            end
        3'h3: // req 1
            begin
            end
        3'h4: // req 1
            begin
            if ((data_chain_combs__taking_transmitter_data!=1'h0))
            begin
                if ((data_transmitter_combs__counter_expired!=1'h0))
                begin
                    data_transmitter_combs__loading_leds__var = 1'h1;
                end //if
            end //if
            end
    //synopsys  translate_off
    //pragma coverage off
        default:
            begin
                if (1)
                begin
                    $display("%t *********CDL ASSERTION FAILURE:led_ws2812_chain:data_transmitter_logic: Full switch statement did not cover all values", $time);
                end
            end
    //pragma coverage on
    //synopsys  translate_on
        endcase
        data_transmitter_combs__idle_transmitter = data_transmitter_combs__idle_transmitter__var;
        data_transmitter_combs__selected_data = data_transmitter_combs__selected_data__var;
        data_transmitter_combs__load_leds = data_transmitter_combs__load_leds__var;
        data_transmitter_combs__drive_bits__valid = data_transmitter_combs__drive_bits__valid__var;
        data_transmitter_combs__drive_bits__value = data_transmitter_combs__drive_bits__value__var;
        data_transmitter_combs__loading_leds = data_transmitter_combs__loading_leds__var;
    end //always

    //b data_transmitter_logic__posedge_clk_active_low_reset_n clock process
        //   
        //       The data transmitter is responsible for reading data bits to the
        //       Neopixel data chain driver (modulator).
        //   
        //       It maintains a shift register (with separate @a red, @a green and @a blue
        //       components), with a @a valid bit.
        //   
        //       Data is loaded into the shift register when it is not valid. The
        //       transmitter then shifts straight in to asking the drive chain to
        //       output @a green[7]. It shifts the @a green bits up every time the
        //       drive chain takes a bit, and after 8 bits it moves to the @a red,
        //       and then the @a blue. At the end of the @a blue it invalidates the
        //       shift register.
        //   
        //       The shift register should be filled quickly enough for the data
        //       chain to not miss a beat, if further LED data is to be driven.
        //   
        //       Instead of driving out a shift register the state machine may be
        //       requested to drive out a 'load leds' value. This is 50us of 'low'
        //       on the output, which is achieved here by roughly 40 sets of drives
        //       of '0' for 1.25us each.
        //       
    always @( posedge clk or negedge reset_n)
    begin : data_transmitter_logic__posedge_clk_active_low_reset_n__code
        if (reset_n==1'b0)
        begin
            data_transmitter_state__shift_register__valid <= 1'h0;
            data_transmitter_state__shift_register__last <= 1'h0;
            data_transmitter_state__shift_register__red <= 8'h0;
            data_transmitter_state__shift_register__green <= 8'h0;
            data_transmitter_state__shift_register__blue <= 8'h0;
            data_transmitter_state__fsm_state <= 3'h0;
            data_transmitter_state__fsm_state <= 3'h0;
            data_transmitter_state__counter <= 6'h0;
        end
        else if (clk__enable)
        begin
            if ((data_transmitter_combs__taking_data!=1'h0))
            begin
                data_transmitter_state__shift_register__valid <= data_state__buffer__valid;
                data_transmitter_state__shift_register__last <= data_state__buffer__last;
                data_transmitter_state__shift_register__red <= data_state__buffer__red;
                data_transmitter_state__shift_register__green <= data_state__buffer__green;
                data_transmitter_state__shift_register__blue <= data_state__buffer__blue;
            end //if
            case (data_transmitter_state__fsm_state) //synopsys parallel_case
            3'h0: // req 1
                begin
                if ((data_state__load_leds!=1'h0))
                begin
                    data_transmitter_state__fsm_state <= 3'h4;
                    data_transmitter_state__counter <= 6'h28;
                end //if
                else
                
                begin
                    if ((data_transmitter_combs__taking_data!=1'h0))
                    begin
                        data_transmitter_state__fsm_state <= 3'h1;
                        data_transmitter_state__counter <= 6'h7;
                    end //if
                end //else
                end
            3'h1: // req 1
                begin
                if ((data_chain_combs__taking_transmitter_data!=1'h0))
                begin
                    data_transmitter_state__counter <= (data_transmitter_state__counter-6'h1);
                    data_transmitter_state__shift_register__green[7:1] <= data_transmitter_state__shift_register__green[6:0];
                    if ((data_transmitter_combs__counter_expired!=1'h0))
                    begin
                        data_transmitter_state__fsm_state <= 3'h2;
                        data_transmitter_state__counter <= 6'h7;
                    end //if
                end //if
                end
            3'h2: // req 1
                begin
                if ((data_chain_combs__taking_transmitter_data!=1'h0))
                begin
                    data_transmitter_state__counter <= (data_transmitter_state__counter-6'h1);
                    data_transmitter_state__shift_register__red[7:1] <= data_transmitter_state__shift_register__red[6:0];
                    if ((data_transmitter_combs__counter_expired!=1'h0))
                    begin
                        data_transmitter_state__fsm_state <= 3'h3;
                        data_transmitter_state__counter <= 6'h7;
                    end //if
                end //if
                end
            3'h3: // req 1
                begin
                if ((data_chain_combs__taking_transmitter_data!=1'h0))
                begin
                    data_transmitter_state__counter <= (data_transmitter_state__counter-6'h1);
                    data_transmitter_state__shift_register__blue[7:1] <= data_transmitter_state__shift_register__blue[6:0];
                    if ((data_transmitter_combs__counter_expired!=1'h0))
                    begin
                        data_transmitter_state__fsm_state <= 3'h0;
                        data_transmitter_state__shift_register__valid <= 1'h0;
                    end //if
                end //if
                end
            3'h4: // req 1
                begin
                if ((data_chain_combs__taking_transmitter_data!=1'h0))
                begin
                    data_transmitter_state__counter <= (data_transmitter_state__counter-6'h1);
                    if ((data_transmitter_combs__counter_expired!=1'h0))
                    begin
                        data_transmitter_state__fsm_state <= 3'h0;
                    end //if
                end //if
                end
    //synopsys  translate_off
    //pragma coverage off
            default:
                begin
                    if (1)
                    begin
                        $display("%t *********CDL ASSERTION FAILURE:led_ws2812_chain:data_transmitter_logic: Full switch statement did not cover all values", $time);
                    end
                end
    //pragma coverage on
    //synopsys  translate_on
            endcase
        end //if
    end //always

    //b data_chain_driver_logic__comb combinatorial process
        //   
        //       The data chain (modulator) starts 'inactive' (it is basically active or
        //       inactive).  It can enter active ONLY on a 400ns clock boundary,
        //       and then only when there is a valid 3-value in hand.  When it
        //       enters 'active' it drives the output pin with @a value[0].
        //   
        //       The data chain is then active for 2 whole 400ns periods; at the
        //       end of the first period it drives out @a value[1], and at the end of
        //       the second period it drives out @a value[2] and becomes inactive, and
        //       invalidates the value-in-hand.
        //   
        //       The value-in-hand can only be loaded if it is invalid - this can
        //       happen during the last 400ns of the previous 'LED data bit'. The
        //       data supplied can be a valid LED 0 or 1 (with the values of 3b100
        //       or 3b110), or it can be part of an LED load train (value of
        //       3b000).
        //       
    always @ ( * )//data_chain_driver_logic__comb
    begin: data_chain_driver_logic__comb_code
        data_chain_combs__clk_enable = (data_chain_state__divider==8'h0);
        data_chain_combs__taking_transmitter_data = (!(data_chain_state__sr__valid!=1'h0)&&(data_transmitter_combs__drive_bits__valid!=1'h0));
        led_chain = data_chain_state__output_data;
    end //always

    //b data_chain_driver_logic__posedge_clk_active_low_reset_n clock process
        //   
        //       The data chain (modulator) starts 'inactive' (it is basically active or
        //       inactive).  It can enter active ONLY on a 400ns clock boundary,
        //       and then only when there is a valid 3-value in hand.  When it
        //       enters 'active' it drives the output pin with @a value[0].
        //   
        //       The data chain is then active for 2 whole 400ns periods; at the
        //       end of the first period it drives out @a value[1], and at the end of
        //       the second period it drives out @a value[2] and becomes inactive, and
        //       invalidates the value-in-hand.
        //   
        //       The value-in-hand can only be loaded if it is invalid - this can
        //       happen during the last 400ns of the previous 'LED data bit'. The
        //       data supplied can be a valid LED 0 or 1 (with the values of 3b100
        //       or 3b110), or it can be part of an LED load train (value of
        //       3b000).
        //       
    always @( posedge clk or negedge reset_n)
    begin : data_chain_driver_logic__posedge_clk_active_low_reset_n__code
        if (reset_n==1'b0)
        begin
            data_chain_state__divider <= 8'h0;
            data_chain_state__output_data <= 1'h0;
            data_chain_state__value_number <= 2'h0;
            data_chain_state__active <= 1'h0;
            data_chain_state__sr__valid <= 1'h0;
            data_chain_state__sr__value <= 3'h0;
        end
        else if (clk__enable)
        begin
            data_chain_state__divider <= (data_chain_state__divider-8'h1);
            if ((data_chain_combs__clk_enable!=1'h0))
            begin
                data_chain_state__divider <= divider_400ns;
            end //if
            if ((data_chain_state__active!=1'h0))
            begin
                if ((data_chain_combs__clk_enable!=1'h0))
                begin
                    data_chain_state__output_data <= data_chain_state__sr__value[data_chain_state__value_number];
                    data_chain_state__value_number <= (data_chain_state__value_number+2'h1);
                    if ((data_chain_state__value_number==2'h2))
                    begin
                        data_chain_state__active <= 1'h0;
                        data_chain_state__sr__valid <= 1'h0;
                    end //if
                end //if
            end //if
            else
            
            begin
                if (((data_chain_state__sr__valid!=1'h0)&&(data_chain_combs__clk_enable!=1'h0)))
                begin
                    data_chain_state__active <= 1'h1;
                    data_chain_state__value_number <= 2'h1;
                    data_chain_state__output_data <= data_chain_state__sr__value[0];
                end //if
            end //else
            if ((!(data_chain_state__sr__valid!=1'h0)&&(data_transmitter_combs__drive_bits__valid!=1'h0)))
            begin
                data_chain_state__sr__valid <= data_transmitter_combs__drive_bits__valid;
                data_chain_state__sr__value <= data_transmitter_combs__drive_bits__value;
            end //if
        end //if
    end //always

endmodule // led_ws2812_chain
